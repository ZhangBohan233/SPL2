/*
 * Superclass of all spl exceptions.
 */
class Exception {
    var message = "";

    /*
     * Create a new <Exception>, with message <msg>.
     */
    fn Exception(msg="") {
        message = msg;
    }
}


/*
 * Exception of assertion failed.
 */
class AssertionException extends Exception {
    fn AssertionException(msg="") {
        Exception(msg);
    }
}


/*
 * Exception of annotations.
 *
 * Exception from all annotations should be derived from this exception.
 */
class AnnotationException extends Exception {
    fn AnnotationException(msg="") {
        Exception(msg);
    }
}


/*
 * A superclass of all iterator classes.
 */
abstract class Iterator {
    abstract fn Iterator();

    abstract fn __more__();

    abstract fn __next__();
}


/*
 * An implementation of a Iterator, works only for integers.
 */
class RangeIterator extends Iterator {

    var iter;
    const step;
    const end;

    /*
     * Creates a new instance.
     *
     * @param begin: the initial value
     * @param end:   the stop value
     * @param step:  the value to be added in each iteration
     */
    fn RangeIterator(begin, end, step) {
        this.iter = begin;
        this.end = end;
        this.step = fn (x) {x + step};
    }

    @Override
    fn __more__() {
        return iter != end;
    }

    @Override
    fn __next__() {
        var temp = iter;
        iter = step(iter);
        return temp;
    }
}


/*
 * Superclass of all iterable classes.
 *
 * Iterable are typically used when calling for (iterable; )
 */
abstract class Iterable {

    /*
     * Returns an object to be iterated, probably an <Iterator>.
     */
    abstract fn __iter__();
}


abstract class OutputStream {
    abstract fn write(obj);

    abstract fn flush();

    abstract fn close();
}

abstract class InputStream {
    abstract fn read();

    abstract fn close();
}

/*
 * Abstract class of lined input stream.
 *
 * All classes extends this must implement <readline>
 */
abstract class LineInputStream extends InputStream {

    /*
     * Returns the next line.
     */
    abstract fn readline();
}

class NativeInputStream extends LineInputStream {

    var ns;

    fn NativeInputStream(stream) {
        ns = stream;
    }

    @Override
    fn readline() {
        return ns.readline();
    }

    @Override
    fn read() {
        return ns.read();
    }

    @Override
    fn close() {
        ns.close();
    }
}

class NativeOutputStream extends OutputStream {

    var ns;

    fn NativeOutputStream(stream) {
        ns = stream;
    }

    @Override
    fn write(obj) {
        ns.write(obj);
    }

    @Override
    fn flush() {
        ns.flush();
    }

    @Override
    fn close() {
        ns.close();
    }
}


class List extends Iterable {

    var arr;
    var length = 0;

    fn List(*args) {
        arr = array(length=8);
        for var x; args {
            append(x);
        }
    }

    fn __getitem__(index) {
        return arr[index];
    }

    fn __setitem__(index, value) {
        arr[index] = value;
    }

    fn __iter__() {
        return to_array();
    }

    fn __str__() {
        return string(to_array());
    }

    fn __repr__() {
        return __str__();
    }

    fn __unpack__() {
        return to_array();
    }

    fn append(v) {
        if length >= arr.size() {
            double_size();
        }
        arr[length] = v;
        length++;
        return this;
    }

    fn insert(index, value) {
        if length >= arr.size() {
            double_size();
        }
        for var i = length + 1; i >= index; i-- {
            arr[i] = arr[i - 1];
        }
        arr[index] = value;
        length++;
    }

    fn pop(index=null) {
        if index === null {
            index = length - 1;
        }
        var val = arr[index];
        for var i = index; i < length; i++ {
            arr[i] = arr[i + 1];
        }
        length--;
        if length < arr.size() / 4 {
            half_size();
        }
        return val;
    }

    fn extend(iter) {
        for var x; iter {
            append(x);
        }
    }

    fn clear() {
        arr = array(length = 8);
    }

    fn copy() {
        return new List(*this);
    }

    fn size() {
        return length;
    }

    /*
     * Swaps the content at index <src> to the content at index <dest>.
     */
    fn swap(src, dest) {
        var temp = this[src];
        this[src] = this[dest];
        this[dest] = temp;
    }

    fn to_array() {
        var s_arr = array(length=length);
        for var i = 0; i < length; i++ {
            s_arr[i] = arr[i];
        }
        return s_arr;
    }

    fn double_size() {
        var big_arr = array(length = arr.size() * 2);
        for var i = 0; i < arr.size(); i++ {
            big_arr[i] = arr[i];
        }
        arr = big_arr;
    }

    fn half_size() {
        var sml_array = array(length = arr.size() / 2);
        for var i = 0; i < sml_arr.size(); i++ {
            sml_arr[i] = arr[i];
        }
        arr = sml_arr;
    }
}


/*
 * Returns a new <List> instance, with initial elements *args
 */
fn list(*args) {
    return new List(*args);
}

/*
 * Returns a <Iterator>, counts from
 */
fn range(n1, n2=null, step=1) {
    var start;
    var stop;
    if n2 === null {
        start = 0;
        stop = n1;
    } else {
        start = n1;
        stop = n2;
    }

}

system.set_in(new NativeInputStream(system.native_in));
system.set_out(new NativeOutputStream(system.native_out));
system.set_err(new NativeOutputStream(system.native_err));
